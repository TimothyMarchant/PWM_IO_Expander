module Main_tb();




endmodule